`timescale 1ns / 1ps

module top_wrapper 
(
    output wire [31:0] o_instruction,
    output wire [15:0] o_process_counter,

    input wire [15:0] i_jmp_address,
    input wire i_en_jmp,

    input wire  i_clk,
    input wire  i_rstn
);


// addi x0, x0, 0        00000000000000000000000000010011
// addi x1, x0, 1        00000000000100000000000010010011
// addi x2, x0, 2        00000000001000000000000100010011
// addi x11, x0, 11      00000000101100000000010110010011
// lw x3, 0(x0)          00000000000000000010000110000011
// sra x4, x3, x11       01000000101100011101001000110011
// beq x4, x1, 30        00000000000100100000111101100011
// sw x3, 0(x1)          00000000001100001010000000100011
// sw x0, 0(x2)          00000000000000010010000000100011
// beq x0, x0, 0         00000000000000000000000001100011
// sw x3, 0(x2)          00000000001100010010000000100011
// sw x0, 0(x1)          00000000000000001010000000100011
// beq x0, x0, 0         00000000000000000000000001100011

localparam MEM_SIZE = 39;
localparam [((32 * MEM_SIZE)-1):0] memory = {
    32'b00000000000000000000000001100011,
    32'b00000000000000000000000000000000,        // nop
    32'b00000000000000000000000000000000,        // nop
    32'b00000000000000001010000000100011,
    32'b00000000000000000000000000000000,        // nop
    32'b00000000000000000000000000000000,        // nop
    32'b00000000001100010010000000100011,
    32'b00000000000000000000000000000000,        // nop
    32'b00000000000000000000000000000000,        // nop
    32'b00000000000000000000000001100011,
    32'b00000000000000000000000000000000,        // nop
    32'b00000000000000000000000000000000,        // nop
    32'b00000000000000010010000000100011,
    32'b00000000000000000000000000000000,        // nop
    32'b00000000000000000000000000000000,        // nop
    32'b00000000001100001010000000100011,
    32'b00000000000000000000000000000000,        // nop
    32'b00000000000000000000000000000000,        // nop
    32'b00000000000100100000111101100011,
    32'b00000000000000000000000000000000,        // nop
    32'b00000000000000000000000000000000,        // nop
    32'b01000000101100011101001000110011,
    32'b00000000000000000000000000000000,        // nop
    32'b00000000000000000000000000000000,        // nop
    32'b00000000000000000010000110000011,
    32'b00000000000000000000000000000000,        // nop
    32'b00000000000000000000000000000000,        // nop
    32'b00000000101100000000010110010011,
    32'b00000000000000000000000000000000,        // nop
    32'b00000000000000000000000000000000,        // nop
    32'b00000000001000000000000100010011,
    32'b00000000000000000000000000000000,        // nop
    32'b00000000000000000000000000000000,        // nop
    32'b00000000000100000000000010010011,
    32'b00000000000000000000000000000000,        // nop
    32'b00000000000000000000000000000000,        // nop
    32'b00000000000000000000000000010011,
    32'b00000000000000000000000000000000,        // nop
    32'b00000000000000000000000000000000         // nop
};

reg [15:0] address = 0;

assign o_process_counter = 0;
assign o_instruction = memory[address+:32];

always @(posedge i_clk) begin
    if (!i_rstn) begin
        address <= 0;
    end else begin
        if (i_en_jmp == 1) begin 
            address <= i_jmp_address << 3;
        end else if (address < (32'h0020 * (MEM_SIZE-1))) begin
            address <= address + 32'h0020; 
        end
    end
end

endmodule
